module top_module ( input a, input b, output out );

    mod_a m0(a,b,out);
	
endmodule